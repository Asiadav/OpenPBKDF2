`define FSB_LEGACY
